`timescale 1ns / 1ps



module skid_buffer#(

    parameter DATAW             = 8,
    parameter PASSTHRU          = 0,
    parameter NOBACKPRESSURE    = 0,
    parameter OUT_REG           = 0

)(
    
    input wire clk,
    input wire reset,
    
    input wire                  valid_in,
    input wire [DATAW-1 : 0]    data_in,
    input wire                  ready_out,
    
    output wire                 ready_in,
    output wire [DATAW-1 : 0]   data_out,
    output wire                 valid_out 
);

    if(PASSTHRU)
    begin
    
        assign valid_out = valid_in;
        assign data_out  = data_in;
        assign ready_in  = ready_out;
            
    end
    else if(NOBACKPRESSURE)
    begin
    
        //The module doesnot use backpressure technique
        //The module doesnot buffer the data , as soon as
        //the input data is valid , the output id produced. 

        
        wire stall = valid_out && ~ready_out;
        
        pipe_register #(
        
            .DATAW  (1 + DATAW),
            .RESETW (1)
            
        ) pipe_reg (
            .clk      (clk),
            .reset    (reset),
            .enable   (!stall),
            .data_in  ({valid_in, data_in}),
            .data_out ({valid_out, data_out})
        );
        
        assign ready_in = ~stall;
    
    end
    else 
    begin
        
        //This module support backpressure which means that if
        //the reciever side cannot handle the requests of the 
        //other side the data will be buffered until the other 
        //side is ready to receive it , this module is usfel for
        //handling the clock domain crossing.
        
        if(OUT_REG)
        begin
            
            reg [DATAW-1 : 0] data_out_r;
            reg [DATAW-1 : 0] buffer;
            reg               valid_out_r;
            reg               use_buffer;
            
            wire push = valid_in && ready_in;
            wire pop  = !valid_out_r || ready_out;
            
            always@(posedge clk)
            begin
            
                if(reset)
                begin
                
                    valid_out_r <= 0;
                    use_buffer  <= 0;
                
                end
                else begin
                
                    if(ready_out)
                    begin
                        
                        //The data is no longer buffered when the other side,
                        //is ready to receive data
                        use_buffer <= 0;
                    
                    end
                    else if(valid_in && valid_out_r)
                    begin
                    
                        //If the receiver on the other side is not ready to receive data,
                        //but there is data available at the input , this data is buffered,
                        //until the receiver on the other side is ready to receive this data.
                        use_buffer <= 1;
                    
                    end
                    
                    if(pop)
                    begin
                    
                        valid_out_r <= valid_in || use_buffer;
                    
                    end
                
                end
            
            end//always end
            
            always@(posedge clk)
            begin
            
                if(push)
                begin
                
                    buffer <= data_in;
                
                end
                if(pop && !use_buffer)
                begin
                
                    data_out_r <= data_in;
                
                end
                else if (ready_out) begin
                        
                    data_out_r <= buffer;  
                
                end
            
            end//always end
            
            assign ready_in  = !use_buffer;
            assign valid_out = valid_out_r;
            assign data_out  = data_out_r;
            
        end//OUT_REG end
        else begin
        
            reg [DATAW-1 : 0] shift_reg [1 : 0];
            reg valid_out_r;
            reg ready_in_r;
            reg rd_ptr_r;
            
            wire push = valid_in && ready_in;
            wire pop  = valid_out_r && ready_out;
            
            always@(posedge clk)
            begin
            
                if(reset)
                begin
                
                    valid_out_r <= 0;
                    ready_in_r  <= 1;
                    rd_ptr_r    <= 1;
                
                end
                else begin
                
                    if(push)
                    begin
                        
                        if(!pop)
                        begin
                            
                            ready_in_r  <= rd_ptr_r;
                            valid_out_r <= 1;     
                        
                        end
                    
                    end//push
                    else if(pop)
                    begin
                    
                        ready_in_r  <= 1;
                        valid_out_r <= rd_ptr_r;
                    
                    end
                    
                    rd_ptr_r <= rd_ptr_r ^ (push ^ pop);
                
                end
            
            end//always end
            
            always @(posedge clk) 
            begin
            
                if (push) 
                begin
                
                    shift_reg[1] <= shift_reg[0];
                    shift_reg[0] <= data_in;
                    
                end
                
            end
            
            assign ready_in  = ready_in_r;
            assign valid_out = valid_out_r;
            assign data_out  = shift_reg[rd_ptr_r];
        
        end
    
    end

endmodule